netcdf idvbad {
dimensions:
	xi_psi = 9 ;
	xi_rho = 10 ;
	xi_u = 9 ;
	xi_v = 10 ;
	eta_psi = 9 ;
	eta_rho = 10 ;
	eta_u = 10 ;
	eta_v = 9 ;
	two = 2 ;
	bath = UNLIMITED ; // (0 currently)
variables:
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	char JPRJ(two) ;
		JPRJ:long_name = "Map projection type" ;
		JPRJ:option\(ME\) = "Mercator" ;
		JPRJ:option\(ST\) = "Stereographic" ;
		JPRJ:option\(LC\) = "Lambert conformal conic" ;
	float PLAT(two) ;
		PLAT:long_name = "Reference latitude(s) for map projection" ;
		PLAT:units = "degree_north" ;
	float PLONG ;
		PLONG:long_name = "Reference longitude for map projection" ;
		PLONG:units = "degree_east" ;
	float ROTA ;
		ROTA:long_name = "Rotation angle for map projection" ;
		ROTA:units = "degree" ;
	char JLTS(two) ;
		JLTS:long_name = "How limits of map are chosen" ;
		JLTS:option\(CO\) = "P1, .. P4 define two opposite corners " ;
		JLTS:option\(MA\) = "Maximum (whole world)" ;
		JLTS:option\(AN\) = "Angles - P1..P4 define angles to edge of domain" ;
		JLTS:option\(LI\) = "Limits - P1..P4 define limits in u,v space" ;
	float P1 ;
		P1:long_name = "Map limit parameter number 1" ;
	float P2 ;
		P2:long_name = "Map limit parameter number 2" ;
	float P3 ;
		P3:long_name = "Map limit parameter number 3" ;
	float P4 ;
		P4:long_name = "Map limit parameter number 4" ;
	float XOFF ;
		XOFF:long_name = "Offset in x direction" ;
		XOFF:units = "meter" ;
	float YOFF ;
		YOFF:long_name = "Offset in y direction" ;
		YOFF:units = "meter" ;
	short depthmin ;
		depthmin:long_name = "Shallow bathymetry clipping depth" ;
		depthmin:units = "meter" ;
	short depthmax ;
		depthmax:long_name = "Deep bathymetry clipping depth" ;
		depthmax:units = "meter" ;
	char spherical ;
		spherical:long_name = "Grid type logical switch" ;
		spherical:option\(T\) = "spherical" ;
		spherical:option\(F\) = "Cartesian" ;
	double hraw(bath, eta_rho, xi_rho) ;
		hraw:long_name = "Working bathymetry at RHO-points" ;
		hraw:units = "meter" ;
		hraw:field = "bath, scalar" ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "Final bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:coordinates = "lon_rho lat_rho" ;
		h:field = "bath, scalar" ;
	double f(eta_rho, xi_rho) ;
		f:long_name = "Coriolis parameter at RHO-points" ;
		f:units = "second-1" ;
		f:field = "Coriolis, scalar" ;
	double pm(eta_rho, xi_rho) ;
		pm:long_name = "curvilinear coordinate metric in XI" ;
		pm:units = "meter-1" ;
		pm:field = "pm, scalar" ;
	double pn(eta_rho, xi_rho) ;
		pn:long_name = "curvilinear coordinate metric in ETA" ;
		pn:units = "meter-1" ;
		pn:field = "pn, scalar" ;
	double dndx(eta_rho, xi_rho) ;
		dndx:long_name = "xi derivative of inverse metric factor pn" ;
		dndx:units = "meter" ;
		dndx:field = "dndx, scalar" ;
	double dmde(eta_rho, xi_rho) ;
		dmde:long_name = "eta derivative of inverse metric factor pm" ;
		dmde:units = "meter" ;
		dmde:field = "dmde, scalar" ;
	double x_rho(eta_rho, xi_rho) ;
		x_rho:long_name = "x location of RHO-points" ;
		x_rho:units = "meter" ;
	double y_rho(eta_rho, xi_rho) ;
		y_rho:long_name = "y location of RHO-points" ;
		y_rho:units = "meter" ;
	double x_psi(eta_psi, xi_psi) ;
		x_psi:long_name = "x location of PSI-points" ;
		x_psi:units = "meter" ;
	double y_psi(eta_psi, xi_psi) ;
		y_psi:long_name = "y location of PSI-points" ;
		y_psi:units = "meter" ;
	double x_u(eta_u, xi_u) ;
		x_u:long_name = "x location of U-points" ;
		x_u:units = "meter" ;
	double y_u(eta_u, xi_u) ;
		y_u:long_name = "y location of U-points" ;
		y_u:units = "meter" ;
	double x_v(eta_v, xi_v) ;
		x_v:long_name = "x location of V-points" ;
		x_v:units = "meter" ;
	double y_v(eta_v, xi_v) ;
		y_v:long_name = "y location of V-points" ;
		y_v:units = "meter" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:option\(0\) = "land" ;
		mask_rho:option\(1\) = "water" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:option\(0\) = "land" ;
		mask_u:option\(1\) = "water" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:option\(0\) = "land" ;
		mask_v:option\(1\) = "water" ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on PSI-points" ;
		mask_psi:option\(0\) = "land" ;
		mask_psi:option\(1\) = "water" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between xi axis and east" ;
		angle:units = "radian" ;

// global attributes:
		:type = "Gridpak file" ;
		:gridid = "                                                                                                                                " ;
		:history = "Created by \"seagrid2roms\" on 01-Mar-2009 12:42:45" ;
		:CPP-options = "DCOMPLEX, DBLEPREC, NCARG_32, PLOTS," ;
data:

 xl = 619188.013259099 ;

 el = 288887.78962873 ;

 JPRJ = "ME" ;

 PLAT = _, _ ;

 PLONG = _ ;

 ROTA = _ ;

 JLTS = "" ;

 P1 = _ ;

 P2 = _ ;

 P3 = _ ;

 P4 = _ ;

 XOFF = _ ;

 YOFF = _ ;

 depthmin = _ ;

 depthmax = _ ;

 spherical = "T" ;

 h =
  190.773685814661, 676.40917538391, 185.589371933765, 179.952627515865, 
    891.531465668186, 1587.25316888552, 3142.45414659357, 3375.24436908043, 
    3745.56151567435, 3969.05080044086,
  753.762224952498, 1207.65474911337, 500.275643069478, 186.2274217176, 
    1005.09712307681, 1707.44378204324, 2642.43517352308, 3350.51821162717, 
    3734.9801743964, 3967.09372980185,
  2008.62916863998, 1595.61059470991, 826.781659657623, 633.888890833158, 
    1108.92300990976, 1607.05027312848, 3150.54031260172, 3339.33217269717, 
    3732.09336517969, 3964.98227017135,
  3294.7083199779, 1994.68670998754, 1091.50429582655, 1006.34851933584, 
    1572.84286486337, 2022.34671229157, 3391.83786094185, 3332.98054334885, 
    3739.85591044992, 3967.51193266832,
  2885.63364048915, 2260.8080008877, 1605.04665769256, 1586.86057606878, 
    1795.08440300572, 2100.06989103826, 3463.62423506393, 3343.65608860733, 
    3746.22272409708, 3971.45575850166,
  3035.43781899047, 2656.00654220132, 2007.90292579215, 1845.79848151114, 
    1996.61054121641, 2259.32835944395, 3513.6714554253, 3307.45167460427, 
    3755.9272005264, 3976.35036508515,
  3078.43994124178, 3430.74108187069, 2279.31179080567, 2023.68629991368, 
    2213.86271286534, 2990.66768074843, 2904.24629617079, 3394.32222566814, 
    3772.3265218775, 3978.95021002981,
  3137.21415453322, 3433.3593203962, 2509.9201534272, 2374.49656724031, 
    2504.08404733515, 3443.62212420656, 3016.94559971624, 3402.378258843, 
    3797.06303613328, 3979.51475262317,
  3192.4513771004, 2952.00782356963, 3512.49895474076, 3401.53944632567, 
    3558.17664935058, 2940.05327984203, 3174.99445644491, 3424.10350458705, 
    3820.81155417451, 3973.78565255103,
  3314.1947158413, 3087.57219479138, 3032.71981888831, 2974.22711397435, 
    3000.15955070688, 3160.59922736022, 3268.71769031304, 3410.28411155159, 
    3805.20636576494, 3964.12249855707 ;

 f =
  1.19643126671356e-05, 1.09025517039847e-05, 9.85578239797317e-06, 
    8.9722245614785e-06, 8.47403064073537e-06, 8.50888410816802e-06, 
    8.93260376563889e-06, 9.53455997827303e-06, 1.01992639495267e-05, 
    1.08511585694005e-05,
  1.22000938731516e-05, 1.11433301403456e-05, 1.01486974038856e-05, 
    9.36942800030595e-06, 8.94549439869812e-06, 8.93857220820034e-06, 
    9.27313516722327e-06, 9.81493458278193e-06, 1.04489535186321e-05, 
    1.11060955274987e-05,
  1.2451681958746e-05, 1.14144330827821e-05, 1.04759442008033e-05, 
    9.78984123177472e-06, 9.42676537034852e-06, 9.38965462758601e-06, 
    9.64823682308626e-06, 1.01290549151857e-05, 1.07300689520009e-05, 
    1.13803248048564e-05,
  1.27088767230481e-05, 1.16999166666459e-05, 1.08172786124264e-05, 
    1.02082323029627e-05, 9.89177307693405e-06, 9.8356600145802e-06, 
    1.00351427570492e-05, 1.04601765962942e-05, 1.10270873591518e-05, 
    1.16626717294276e-05,
  1.29701020397239e-05, 1.19959495857903e-05, 1.11668956922621e-05, 
    1.06212632709955e-05, 1.03410886140052e-05, 1.02740755141339e-05, 
    1.04287489095966e-05, 1.08047993174011e-05, 1.13371732535447e-05, 
    1.1951574227218e-05,
  1.32346317507431e-05, 1.2299887043752e-05, 1.15207734428595e-05, 
    1.10270267988992e-05, 1.07756300210746e-05, 1.07038169406954e-05, 
    1.08259179148857e-05, 1.11606513872509e-05, 1.16587747515307e-05, 
    1.22459304134759e-05,
  1.35030096176825e-05, 1.26110151217239e-05, 1.18772533737824e-05, 
    1.14259665401288e-05, 1.11981643772647e-05, 1.11262870652723e-05, 
    1.12261991660486e-05, 1.15275465142112e-05, 1.1992271219544e-05, 
    1.25461596871091e-05,
  1.37780795160719e-05, 1.29317564376177e-05, 1.22374954792137e-05, 
    1.18207990489298e-05, 1.16131248148713e-05, 1.15454450637333e-05, 
    1.16325698369259e-05, 1.19087271276092e-05, 1.23415471973498e-05, 
    1.28546052304926e-05,
  1.40627134274682e-05, 1.32642332516607e-05, 1.26019863037975e-05, 
    1.22129540855737e-05, 1.20231601578589e-05, 1.19639663661421e-05, 
    1.20472989815203e-05, 1.23068608407691e-05, 1.27099708013758e-05, 
    1.31733396699348e-05,
  1.4383724778419e-05, 1.36413952312666e-05, 1.29968117041988e-05, 
    1.26293330713952e-05, 1.24568340710612e-05, 1.2413727163731e-05, 
    1.2505422935536e-05, 1.27588792295629e-05, 1.31367864801847e-05, 
    1.35265517152389e-05 ;

 pm =
  1.45578461805502e-05, 1.42881683468219e-05, 1.44641276001386e-05, 
    1.47720244298872e-05, 1.50217011035432e-05, 1.47036675110423e-05, 
    1.44604949950046e-05, 1.43187920218189e-05, 1.42605943621137e-05, 
    1.44937814596955e-05,
  1.51020785017955e-05, 1.43735907521456e-05, 1.49242212955364e-05, 
    1.58958762457195e-05, 1.65725233791168e-05, 1.57527284126229e-05, 
    1.49055278083044e-05, 1.44587980540838e-05, 1.42630550569951e-05, 
    1.49325574752812e-05,
  1.56531804570391e-05, 1.45844839300233e-05, 1.55089402266866e-05, 
    1.71465227849946e-05, 1.82370076263428e-05, 1.69243954059851e-05, 
    1.54576278393595e-05, 1.46639161092297e-05, 1.43357130651605e-05, 
    1.53784377986342e-05,
  1.62425867087434e-05, 1.49118209581042e-05, 1.61949201270547e-05, 
    1.84622788690832e-05, 1.99225906219439e-05, 1.81569156362851e-05, 
    1.60877049309362e-05, 1.49280750088227e-05, 1.44759413503257e-05, 
    1.58491032159376e-05,
  1.68938397827088e-05, 1.53421497380487e-05, 1.6975612828717e-05, 
    1.98391615773246e-05, 2.16267128695056e-05, 1.94407450333828e-05, 
    1.67837617657411e-05, 1.52449573286819e-05, 1.46746239338919e-05, 
    1.63651616165459e-05,
  1.76325169890752e-05, 1.58622211038046e-05, 1.78509448342348e-05, 
    2.12919525081461e-05, 2.33742681352902e-05, 2.07826478745288e-05, 
    1.75396600528617e-05, 1.56067555023573e-05, 1.49204434038738e-05, 
    1.69516954551355e-05,
  1.8492901368266e-05, 1.64569430904834e-05, 1.88274622235018e-05, 
    2.28524823946171e-05, 2.52107129887131e-05, 2.22030532242131e-05, 
    1.83537261119933e-05, 1.6003931835486e-05, 1.51985959762476e-05, 
    1.76448066021387e-05,
  1.95294131273276e-05, 1.71030415026329e-05, 1.99216120729193e-05, 
    2.45776487470717e-05, 2.72096217801843e-05, 2.37404599629798e-05, 
    1.92289258978696e-05, 1.64244959737476e-05, 1.54864602415611e-05, 
    1.85011740691429e-05,
  2.08415690740406e-05, 1.77544488770923e-05, 2.11723330454648e-05, 
    2.65780660070051e-05, 2.95056417208437e-05, 2.54695564006318e-05, 
    2.01766106480044e-05, 1.68534077487494e-05, 1.57438504217612e-05, 
    1.96203040973059e-05,
  2.26182069759159e-05, 1.83007860510638e-05, 2.27458205150673e-05, 
    2.92213345837385e-05, 3.25300817004873e-05, 2.76440881766263e-05, 
    2.12656539736031e-05, 1.72830324096374e-05, 1.58787701611721e-05, 
    2.11776010096472e-05 ;

 pn =
  6.94749276209715e-05, 7.81414667526562e-05, 6.76020395263691e-05, 
    5.61654375911629e-05, 5.18359138022938e-05, 5.71228990815996e-05, 
    6.92610999667815e-05, 8.23158424356185e-05, 9.13934051762509e-05, 
    8.13531612890682e-05,
  6.42285477978207e-05, 6.60118281188647e-05, 5.8556438021378e-05, 
    5.05996099685718e-05, 4.75984245669992e-05, 5.1289064325796e-05, 
    5.99152739585199e-05, 6.96900442073516e-05, 7.67088968227649e-05, 
    7.41856504991729e-05,
  6.2347388168969e-05, 6.23579629017425e-05, 5.65626480313114e-05, 
    5.05643780934262e-05, 4.83267184489287e-05, 5.10932130253728e-05, 
    5.7744115870858e-05, 6.56858453118895e-05, 7.17424755425562e-05, 
    7.17302705395132e-05,
  6.1330845870713e-05, 6.05641652127262e-05, 5.60030371104035e-05, 
    5.14719043306592e-05, 4.98014726684056e-05, 5.18525870923785e-05, 
    5.69769839810821e-05, 6.34389516468291e-05, 6.88053392820823e-05, 
    7.00666626533854e-05,
  6.07015511513837e-05, 5.95478601272663e-05, 5.59909148902241e-05, 
    5.2635083723553e-05, 5.13983491545106e-05, 5.28537184749713e-05, 
    5.66961807861711e-05, 6.18598122903361e-05, 6.66734024999018e-05, 
    6.8883452929879e-05,
  6.02217724387054e-05, 5.8818969865999e-05, 5.61332321021063e-05, 
    5.37694054355552e-05, 5.28666315235748e-05, 5.37924001337667e-05, 
    5.64930945527035e-05, 6.04626754995072e-05, 6.48070937635371e-05, 
    6.7818453507346e-05,
  5.97087171671768e-05, 5.80275621133835e-05, 5.61540809483614e-05, 
    5.46866129122834e-05, 5.40449018371329e-05, 5.44595541142509e-05, 
    5.60812019701418e-05, 5.89074367082835e-05, 6.28366414016225e-05, 
    6.67158663593564e-05,
  5.89218426453559e-05, 5.67485051587649e-05, 5.57145636856738e-05, 
    5.51417682878712e-05, 5.47140061049007e-05, 5.45817364448286e-05, 
    5.51131488192071e-05, 5.67973187324563e-05, 6.03302141686888e-05, 
    6.53816723199753e-05,
  5.7316240287628e-05, 5.40979467569047e-05, 5.40674019582471e-05, 
    5.45085041009504e-05, 5.42765023545189e-05, 5.34882139015041e-05, 
    5.28403752580477e-05, 5.33357497639084e-05, 5.64084306849541e-05, 
    6.32627963253437e-05,
  5.14662491795904e-05, 4.50146141051879e-05, 4.63681823269544e-05, 
    4.80525820981648e-05, 4.80444156871333e-05, 4.64437854516509e-05, 
    4.45367936708363e-05, 4.37867208555247e-05, 4.59645200057035e-05, 
    5.69133343509269e-05 ;

 dndx =
  0, 199.385665253394, 2503.62062874801, 2249.59548729033, -149.214810748625, 
    -2426.76256799867, -2678.89225604782, -1748.20521600389, 
    71.8777725146892, 0,
  0, 754.070373548739, 2307.09895498998, 1965.77860666401, -132.832265415411, 
    -2159.4318737338, -2574.04087201878, -1826.96872870258, 
    -434.778065155934, 0,
  0, 820.173740943939, 1870.16209084628, 1506.48769901264, -102.34868200275, 
    -1687.35266011261, -2174.04553329415, -1689.51891323281, 
    -641.432191152856, 0,
  0, 775.582671934495, 1458.33037229353, 1111.77652551786, -71.3169152157388, 
    -1264.39047597855, -1761.12736885381, -1508.59536293724, 
    -745.531740585629, 0,
  0, 692.998384491528, 1102.76008038096, 797.918714968295, -39.2950940183528, 
    -909.002717407697, -1377.28026975433, -1319.69388462972, 
    -824.154777712344, 0,
  0, 604.734448010831, 798.309456772298, 550.382162382299, -3.97504053798184, 
    -607.122396474821, -1025.42873708539, -1135.43446351798, 
    -896.939964859361, 0,
  0, 530.085716170017, 526.410478874033, 347.494079652763, 38.1200298471904, 
    -335.923006410774, -693.232815847667, -958.502680182186, 
    -993.423549506503, 0,
  0, 488.496758030553, 256.7317902086, 164.113702207702, 93.0367837850499, 
    -66.1826985992375, -357.340883348514, -784.523919614978, 
    -1155.8294164465, 0,
  0, 524.185385523058, -69.6143518125391, -35.6268565725368, 
    174.973129553366, 250.371640043832, 26.7215228830046, -598.537941601189, 
    -1471.03590840291, 0,
  0, 1068.15171147871, -702.235753832145, -376.219668669064, 
    360.434884344586, 819.6358166523, 653.284094212691, -348.717142779156, 
    -2633.69967161678, 0 ;

 dmde =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -2403.34968256894, -710.979160130286, -2328.80996166322, -4687.33290589028, 
    -5868.39974949644, -4461.96865784413, -2230.47325215714, 
    -821.843126220716, -183.721997615714, -1984.49801602079,
  -2324.75131363521, -1255.57342633868, -2628.7067744616, -4372.45164452573, 
    -5073.28286368428, -4202.81649409776, -2464.96696742285, 
    -1087.08431896704, -515.535208905283, -1936.35623873307,
  -2345.80326034186, -1693.05243915508, -2785.4514935393, -3957.75336874174, 
    -4297.22254390358, -3823.97390033962, -2555.79041311705, 
    -1299.57325919677, -805.506818100861, -1960.34765196646,
  -2426.57386537426, -2009.0087058922, -2864.15685296026, -3599.19650052051, 
    -3706.09361182659, -3479.1847072112, -2572.8112938798, -1456.52832927982, 
    -1028.99966059729, -2051.95154189921,
  -2559.18552192661, -2207.64374050333, -2897.06621769287, -3323.21683054368, 
    -3286.71750045447, -3199.75356072856, -2548.27469235357, 
    -1555.40785160362, -1174.64779693955, -2215.75787925944,
  -2754.29245948814, -2286.87054132193, -2911.35141259839, -3139.36341587519, 
    -3015.19144734414, -2997.44053159266, -2504.33145261795, 
    -1595.07393700404, -1224.800805846, -2470.26280993353,
  -3046.88536779163, -2220.35769831366, -2941.2261944505, -3066.95610459989, 
    -2886.92680741559, -2888.14509899674, -2461.25553094407, 
    -1574.73199789643, -1139.34380204593, -2853.14504782232,
  -3496.32311558287, -1913.33543062114, -3116.31007969485, -3232.90136463323, 
    -3005.46393732187, -2974.041702558, -2490.40102066734, -1512.22613717467, 
    -797.682876563511, -3415.46112093202,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 x_rho =
  -5583428.39066481, -5531345.89610071, -5478506.38581839, -5421685.23845359, 
    -5358335.72997491, -5291131.95036392, -5224632.62729462, 
    -5160058.97434061, -5096024.10836984, -5032118.14800688,
  -5573426.06539198, -5522319.55660065, -5468818.98143168, -5413320.24541145, 
    -5355067.90480094, -5293571.02084097, -5229513.5620912, 
    -5165275.11533243, -5100805.35224214, -5037664.44552498,
  -5562560.85344831, -5512370.07704856, -5458895.55763871, -5405244.54440801, 
    -5351693.80008721, -5295388.18311458, -5234161.97765047, 
    -5170679.15145662, -5106115.6268986, -5043749.26746132,
  -5551293.21653312, -5502156.91904634, -5449325.93578584, -5397853.24116121, 
    -5348405.31740076, -5296564.21540613, -5238283.13680194, 
    -5175929.93799002, -5111606.04990786, -5050107.12232544,
  -5539774.73515905, -5491836.63135547, -5440131.45903534, -5391034.41953517, 
    -5345214.23812032, -5297262.93304832, -5241924.74277605, 
    -5180989.22473518, -5117179.55328244, -5056642.53699884,
  -5528116.38478599, -5481508.86408877, -5431294.90716158, -5384693.17070336, 
    -5342129.76561966, -5297617.76080036, -5245158.27290443, 
    -5185849.31992841, -5122761.3717232, -5063263.34752767,
  -5516380.49341508, -5471195.24124214, -5422737.68016338, -5378717.59766579, 
    -5339149.52319524, -5297751.8435135, -5248088.71514717, 
    -5190546.58415452, -5128308.04584474, -5069900.36977858,
  -5504575.10810872, -5460820.1677548, -5414315.53235764, -5372986.25394197, 
    -5336265.32508489, -5297779.46541917, -5250849.05888412, 
    -5195166.4919484, -5133809.07394201, -5076480.29213617,
  -5492732.417041, -5450320.06105164, -5405896.28353273, -5367409.41485196, 
    -5333484.46927464, -5297810.17564897, -5253572.08548357, 
    -5199798.57791817, -5139234.63210693, -5082899.66298808,
  -5480361.13007459, -5438726.67152955, -5396647.21165659, -5361534.46236217, 
    -5330687.19224091, -5298045.64249925, -5256683.59522753, 
    -5204959.1488041, -5144892.48484172, -5089099.45731772 ;

 y_rho =
  524556.30099717, 477822.625077906, 431798.244355935, 392985.26404336, 
    371113.353120532, 372643.334707119, 391245.44459485, 417684.045288262, 
    446895.249677081, 475561.666791859,
  534941.802844045, 488416.036467306, 444672.394673554, 410429.900064051, 
    391811.480081184, 391507.560886528, 406200.288223113, 430003.25926074, 
    457872.945380064, 486777.47773017,
  546026.602030676, 500346.834250716, 459059.698735102, 428900.522830504, 
    412948.527035973, 411318.340890469, 422678.427990539, 443808.97722074, 
    470235.517244142, 498845.337002758,
  557361.862810003, 512914.285599011, 474071.349567965, 447289.489864738, 
    433379.93783867, 430913.988529742, 439681.055213512, 458366.427629731, 
    483301.301565556, 511274.161332185,
  568878.380873779, 525950.316540545, 489452.703430319, 465450.148942351, 
    453130.280576906, 450184.073448215, 456984.521683614, 473522.499691826, 
    496946.236541438, 523995.571773702,
  580544.37702758, 539338.987336798, 505027.306782478, 483298.610112842, 
    472239.462209526, 469080.871144105, 474451.434544469, 489178.037181052, 
    511102.702202374, 536961.418647825,
  592384.044523856, 553049.310372306, 520722.512781383, 500854.268520897, 
    490828.732407894, 487665.934540961, 492062.40038588, 505325.563345994, 
    525788.065098194, 550190.527406131,
  604523.167379377, 567188.628428304, 536589.7799136, 518236.667507357, 
    509092.916654609, 506113.491120649, 509948.976409376, 522108.699307283, 
    541174.272804577, 563786.612265104,
  617088.867522802, 581851.102793379, 552650.868665139, 535508.736040319, 
    527148.445765065, 524541.383280222, 528211.625203389, 539645.886035975, 
    557410.688769066, 577841.540895123,
  631266.254205807, 598491.946410402, 570056.654013016, 553856.482589712, 
    546254.228827995, 544354.73382056, 548395.46815758, 559566.745520553, 
    576229.750555463, 593423.448109016 ;

 x_psi =
  -5553079.49266222, -5500567.40303947, -5446221.22578351, -5387665.2837307, 
    -5324912.48945707, -5259665.67348953, -5194711.96837775, 
    -5130520.22119864, -5066267.46824602,
  -5543404.08386573, -5490691.43148305, -5436705.06401741, -5381401.01868419, 
    -5324588.87158017, -5263543.73570332, -5199976.8133717, 
    -5135822.17704062, -5071443.93105514,
  -5533059.35848983, -5480671.10625543, -5427654.75933826, -5375626.91777676, 
    -5323805.30832777, -5266776.57348701, -5205008.2009387, 
    -5141237.63889425, -5077035.62858357,
  -5522364.44870329, -5470741.39016891, -5419175.6273978, -5370320.68101791, 
    -5322706.99315409, -5269402.2555435, -5209703.03783289, 
    -5146630.96270753, -5082860.02066417,
  -5511489.46428832, -5460976.53999409, -5411219.87472605, -5365399.5251229, 
    -5321410.40740004, -5271533.00006309, -5214064.14062849, 
    -5151948.33560045, -5088801.28599685,
  -5500522.739771, -5451371.04998623, -5403690.86288319, -5360781.01422607, 
    -5320003.28491031, -5273296.54068671, -5218143.63604149, 
    -5157177.05962134, -5094774.95020022,
  -5489493.43205066, -5441860.30877033, -5396471.13533532, -5356392.84871503, 
    -5318554.64620678, -5274823.29961494, -5222026.15407999, 
    -5162335.10493048, -5100710.01232789,
  -5478363.23904171, -5432302.42844619, -5389414.65760013, -5352165.59450535, 
    -5317125.12178147, -5276253.77177775, -5225834.44050813, -5167479.492265, 
    -5106538.63352032,
  -5466940.11040557, -5422372.42794294, -5382282.45821146, -5348001.62120731, 
    -5315775.63190987, -5277771.97067818, -5229775.52747798, 
    -5172757.74209878, -5112201.26639824 ;

 y_psi =
  506402.439237972, 459794.172183729, 418195.955160872, 388813.161775744, 
    378990.550537557, 388681.610123952, 410269.903865647, 437708.302378139, 
    466615.514280336,
  517388.240071274, 472102.786970363, 434054.877075615, 409021.536035844, 
    399975.807622937, 406385.842217417, 424700.654728536, 450052.007331468, 
    478250.304701161,
  529048.073830635, 485362.163836719, 450613.006308245, 429021.791594622, 
    420661.97367347, 424670.516858956, 440080.389122809, 463366.289182256, 
    490659.193223733,
  541117.861965085, 499209.907633539, 467404.506545222, 448496.05078399, 
    440744.772501805, 443073.313461592, 456039.345926244, 477371.19069386, 
    503582.994654018,
  553488.694166482, 513450.336604957, 484215.461083613, 467408.979338281, 
    460212.311169943, 461416.071594347, 472407.845751533, 491948.297586904, 
    516924.482673104,
  566136.794503714, 527984.793326526, 500960.156017364, 485823.398608835, 
    479152.235313685, 479660.903411632, 489127.503164079, 507072.138896499, 
    530674.852479626,
  579116.607892048, 542795.628935965, 517638.021022665, 503849.174460585, 
    497700.594923879, 497864.942627906, 506233.011425099, 522803.470272341, 
    544903.253879225,
  592606.175419366, 557969.838508196, 534339.79561217, 521653.408389791, 
    516056.67704665, 516196.056132184, 523885.586371227, 539332.937307985, 
    559798.947765757,
  607095.852712689, 573832.443447021, 551363.349562975, 539580.956412646, 
    534618.232170309, 535084.226880557, 542546.956520637, 557169.860743101, 
    575858.815634912 ;

 x_u =
  -5557371.4938387, -5505148.70696928, -5450862.79144424, -5390817.46527348, 
    -5324869.9453845, -5257607.63315946, -5192167.49801711, 
    -5128073.50861833, -5063990.27844043,
  -5548376.05233146, -5495698.12824881, -5441451.98673086, -5384497.12504679, 
    -5324815.24389277, -5261666.61130871, -5197344.60736729, 
    -5133129.8028649, -5068776.95865555,
  -5538285.64226975, -5485673.25396372, -5432102.52647501, -5378446.22373083, 
    -5324245.77416575, -5265244.94487507, -5202535.31989816, 
    -5138530.0974343, -5074204.13948272,
  -5527744.26803246, -5475689.75104548, -5423347.00616435, -5372921.54294869, 
    -5323287.36200593, -5268157.98924234, -5207397.90495881, 
    -5143940.67619894, -5079926.15348862,
  -5516942.42479986, -5465837.16550899, -5415137.42807671, -5367817.01898496, 
    -5322077.55444341, -5270521.82358908, -5211922.99098496, 
    -5149300.74145516, -5085821.89028156,
  -5506013.79490156, -5456155.90566741, -5407408.55291256, -5363056.96526664, 
    -5320716.02096833, -5272452.71554199, -5216134.74880032, 
    -5154573.6779303, -5091788.86438356,
  -5495019.71735869, -5446613.7453822, -5400052.57624126, -5358563.36179337, 
    -5319280.43199565, -5274080.43829343, -5220101.52072905, 
    -5159760.81654103, -5097750.5853748,
  -5483935.41756721, -5437089.14028394, -5392926.20354139, -5354260.08346909, 
    -5317833.24415842, -5275543.41863165, -5223934.63752482, 
    -5164909.00747523, -5103645.5513252,
  -5472759.3980351, -5427465.49772071, -5385910.92941942, -5350099.65801804, 
    -5316438.28893944, -5276976.03135457, -5227749.03405246, 
    -5170061.97071006, -5109379.09321282,
  -5460680.02058561, -5416774.48779129, -5378369.93501455, -5345798.09902477, 
    -5315138.75607383, -5278713.38831833, -5232029.43967928, 
    -5175689.57768902, -5115050.61449612 ;

 y_u =
  501471.773765126, 454345.861562779, 411015.552629259, 379222.632178042, 
    368997.117068537, 380586.304560291, 403815.762709774, 432228.602718235, 
    461408.293995344,
  511758.961870284, 465769.898689811, 425955.266878506, 398846.351863028, 
    389420.67034244, 397370.272598262, 417298.055304111, 443703.572220739, 
    472282.459499295,
  523161.599376964, 478647.974342785, 442292.732073926, 419091.369211735, 
    410400.232831761, 415504.195844601, 432309.319939051, 456617.144731159, 
    484385.949681669,
  535039.080740229, 492225.447486568, 458994.027267651, 438826.389797589, 
    430778.934937608, 433869.341816102, 447998.822236289, 470290.387965578, 
    497063.361924892,
  547268.759854536, 506289.081634851, 475815.30057909, 458020.682858185, 
    450551.937520832, 452257.188289039, 464178.19194183, 484591.596165158, 
    510203.741189081,
  559777.837261677, 520684.797805109, 492598.822639591, 476673.489146632, 
    469741.706658735, 470550.314597388, 480725.072605859, 499441.559690829, 
    523747.426347182,
  572572.479757712, 535348.417768914, 509299.623973841, 494871.600308817, 
    488459.977912871, 488755.138474785, 497619.690436034, 514847.752582082, 
    537715.423052946,
  585797.634293519, 550342.767013041, 525991.847542102, 512781.555658691, 
    506903.892149852, 507017.454832962, 514994.324109234, 530969.960703119, 
    552268.366027587,
  599594.065990577, 565708.387677577, 542709.646880446, 530497.647128935, 
    525197.918838491, 525443.55491515, 532953.289252055, 547944.826353829, 
    567546.651080343,
  615516.760287374, 582676.655909788, 560621.393517919, 549228.463292815, 
    544671.143042216, 545512.714554385, 553091.870127881, 567450.225037136, 
    585156.703012269 ;

 x_v =
  -5578583.23717002, -5527021.29293238, -5473765.78964038, -5417525.9534213, 
    -5356739.09808985, -5292414.6145433, -5227061.81872203, 
    -5162602.91976899, -5098310.68995105, -5034795.27953722,
  -5568056.70248407, -5517392.86370256, -5463819.87359425, -5409193.20430302, 
    -5353372.3348437, -5294569.49079731, -5231903.17691409, 
    -5167990.76121461, -5103429.33400769, -5040666.02356761,
  -5556967.73468123, -5507286.80430273, -5454065.84151042, -5401472.47777078, 
    -5350038.62093506, -5296044.60514266, -5236285.25855124, 
    -5173325.95552905, -5108844.2341111, -5046898.93579742,
  -5545556.27377484, -5497000.61367575, -5444679.94513115, -5394376.67251909, 
    -5346796.29940304, -5296964.92848092, -5240161.04153519, 
    -5178485.86831814, -5114388.5212719, -5053359.75663274,
  -5533958.74094516, -5486671.59950737, -5435673.11218882, -5387811.76773415, 
    -5343658.95986457, -5297475.05815968, -5243586.06217214, 
    -5183442.3155151, -5119972.33068315, -5059946.40063398,
  -5522255.26240122, -5476350.76094144, -5426987.27284024, -5381666.11644681, 
    -5340626.69992373, -5297705.3693216, -5246654.40266476, -5188215.0711794, 
    -5125541.24900916, -5066584.38985576,
  -5510487.79100315, -5466023.7276231, -5418521.34196055, -5375829.59143415, 
    -5337696.11581974, -5297771.79755588, -5249480.66354358, 
    -5192858.9465349, -5131063.83396478, -5073202.43720793,
  -5498658.76319459, -5455595.13800529, -5410118.02877487, -5370185.4734718, 
    -5334861.74591965, -5297786.90584645, -5252204.95405399, 
    -5197472.4650153, -5136531.79326983, -5079717.5271265,
  -5486680.73417834, -5444783.11610959, -5401475.94525861, -5364563.61700151, 
    -5332104.82254593, -5297883.49913786, -5255032.68192891, 
    -5202251.50209653, -5141991.11435271, -5086026.04094327 ;

 y_v =
  529609.186262504, 482873.876575468, 437950.490135666, 401447.729124311, 
    381257.894900019, 381816.059836955, 398420.710859171, 423574.05606092, 
    452132.548398569, 481003.123825779,
  540444.791232427, 494286.248348935, 451765.26911692, 419657.181328962, 
    402460.517586842, 401423.201254296, 414351.69453254, 436797.17620446, 
    463953.022436953, 492759.48951755,
  551666.926291372, 506560.8299424, 466503.365285522, 438113.056260438, 
    423247.470832239, 421148.32595227, 431127.908229086, 451002.428685928, 
    476687.790914601, 505016.865209912,
  563101.900904134, 519384.595277297, 481731.232063587, 456408.65632593, 
    443342.579971097, 440598.118237193, 448308.868813676, 465879.79764759, 
    490059.271893216, 517604.61402968,
  574691.656426668, 532603.317096491, 497221.395351804, 474412.479039027, 
    462756.785676896, 459675.530049279, 465699.797709547, 481289.117576543, 
    503960.213365718, 530446.920813435,
  586439.361761783, 546153.498244394, 512861.964734238, 492110.396321407, 
    481591.298110483, 478406.99119253, 483237.373676298, 497188.229783719, 
    518375.647599394, 543540.769996979,
  598404.148825127, 560053.26196269, 528627.03269036, 509556.073701011, 
    499986.387502422, 496891.833725959, 500957.471290837, 513622.90716261, 
    533376.809502253, 556932.687499868,
  610737.380093442, 574440.056175187, 544588.766455334, 526877.524075672, 
    518134.913191969, 515316.300254264, 519018.868025251, 530766.65163637, 
    549167.156494246, 570744.681058726,
  623830.125624462, 589739.599615638, 561034.663722179, 544394.251540049, 
    536409.544249702, 534096.185692581, 537866.271867875, 549101.89072853, 
    566279.895165685, 585307.892048735 ;

 lat_rho =
  4.70697053176975, 4.28843502205269, 3.87603348787565, 3.52809061090347, 
    3.33196133176428, 3.34568116728333, 3.5124911876455, 3.74952101323725, 
    4.01133361247221, 4.2681823611482,
  4.79994649162288, 4.38332656052886, 3.99141365827055, 3.68449144806798, 
    3.51756643414371, 3.51484105462397, 3.64657318414857, 3.85994466241495, 
    4.10970234871004, 4.36865150173907,
  4.89916958203408, 4.4901835151592, 4.12033643118514, 3.85006123620059, 
    3.70707056711782, 3.69245650931878, 3.79429016850242, 3.98367591636756, 
    4.22046628670085, 4.47673866683453,
  5.00061910335757, 4.60272561837611, 4.25483146786859, 4.01486661532993, 
    3.89020947524026, 3.86810779902115, 3.94668221628759, 4.11412412164902, 
    4.33751342726123, 4.58804208023829,
  5.10367455426639, 4.71944523879549, 4.3926144616106, 4.17759327162267, 
    4.06720597266926, 4.04080543029565, 4.10174200995566, 4.24991387724661, 
    4.45972948228247, 4.70194771937913,
  5.20805048954048, 4.8393018855289, 4.53210249963857, 4.33748956022691, 
    4.23841954748527, 4.21012191548948, 4.25823588952745, 4.39015337974632, 
    4.58650574329523, 4.81802274722185,
  5.31396251416008, 4.96201612240547, 4.67264346200181, 4.49472984539672, 
    4.40493858042502, 4.37660943797113, 4.41598827746869, 4.53477250192608, 
    4.71799481608375, 4.93643416565447,
  5.42253437000458, 5.0885458826332, 4.814696281516, 4.650384686497, 
    4.56850904736286, 4.54182830976944, 4.57617485479382, 4.68505322040592, 
    4.85573206020886, 5.05810812893291,
  5.53490177167642, 5.21973147565454, 4.95845468338179, 4.80501804079035, 
    4.73017477893198, 4.70683398357099, 4.73969322136479, 4.84205222449025, 
    5.001050691845, 5.18386483969784,
  5.66165586207369, 5.36858178821929, 5.11421265517549, 4.96924174093514, 
    4.90120166144818, 4.8841997652097, 4.92036622798026, 5.02034422172025, 
    5.16944151458889, 5.32325397695204 ;

 lon_rho =
  -50.1578679834768, -49.6899929246753, -49.215317331901, -48.704873316364, 
    -48.1357827754333, -47.5320679841136, -46.934681569509, -46.354594115447, 
    -45.7793467711681, -45.2052574305397,
  -50.0680136367458, -49.6089061956371, -49.1282920283896, -48.6297276912511, 
    -48.1064267718813, -47.5539789976397, -46.9785286946145, 
    -46.4014525137187, -45.8222983382277, -45.2550817390551,
  -49.9704076806644, -49.5195265802896, -49.0391464809364, -48.5571808765589, 
    -48.076116022472, -47.5703031947185, -47.020287019006, -46.4499988389386, 
    -45.8700023717601, -45.3097437986413,
  -49.8691866019052, -49.4277782502445, -48.9531792586558, -48.4907822435794, 
    -48.0465744453419, -47.5808678994656, -47.0573088167609, 
    -46.4971684700907, -45.9193247402412, -45.3668586074325,
  -49.7657121006298, -49.3350675371608, -48.870582094555, -48.4295264109635, 
    -48.0179078766902, -47.587144721662, -47.0900226224941, 
    -46.5426177924243, -45.9693934483731, -45.4255684973908,
  -49.6609811077698, -49.242289632461, -48.7912002933924, -48.3725607799028, 
    -47.9901989936058, -47.5903322620581, -47.1190705417924, 
    -46.5862777081665, -46.0195368536199, -45.4850455278483,
  -49.5555535373125, -49.1496387919779, -48.7143277641776, -48.3188801409525, 
    -47.9634264453391, -47.591536773436, -47.1453957178062, 
    -46.6284748570242, -46.0693645452942, -45.5446681938113,
  -49.4495016788019, -49.0564359191396, -48.638668698059, -48.2673934983821, 
    -47.9375166963579, -47.5917849105663, -47.1701928401224, 
    -46.6699770863012, -46.1187821829481, -45.6037779116873,
  -49.3431146897367, -48.9621098296871, -48.5630356744877, -48.217294824365, 
    -47.9125353069942, -47.5920607911802, -47.1946547296881, 
    -46.7115887163435, -46.1675218481021, -45.6614453398691,
  -49.2319791409251, -48.8579624026148, -48.4799480634943, -48.16451809459, 
    -47.8874064001015, -47.5941760713208, -47.2226064976785, 
    -46.7579479091377, -46.2183482957048, -45.7171402362219 ;

 lat_psi =
  4.54441599467746, 4.12691695157124, 3.75410987699649, 3.4906816723302, 
    3.40260137433856, 3.48950209013985, 3.68305732913646, 3.92900212711403, 
    4.18803417284481,
  4.64278822333717, 4.23719506301298, 3.89625863952433, 3.67186590077906, 
    3.59076815211154, 3.64823684498754, 3.81241649983544, 4.0396218765728, 
    4.29226742508688,
  4.74718106358124, 4.35597385238667, 4.04464898815573, 3.8511479896052, 
    3.77621515822493, 3.8121463600117, 3.95026104853765, 4.15892266159351, 
    4.40341994345005,
  4.85522766812053, 4.48000326160114, 4.19510300507859, 4.02567878774903, 
    3.95621523329186, 3.97708321223532, 4.09327279950328, 4.28439214960744, 
    4.51916713366256,
  4.96595120525286, 4.6075278734124, 4.34570231098279, 4.19514307806963, 
    4.13066349009954, 4.14144912269912, 4.23992801629744, 4.41496614048369, 
    4.63863578821256,
  5.07913717337621, 4.73766194829325, 4.49567814043682, 4.36010530381038, 
    4.30034701175143, 4.30490367481874, 4.38970073191983, 4.55041319985606, 
    4.76174469292531,
  5.19527092997449, 4.87024537950666, 4.64502472566484, 4.52155088086932, 
    4.4664858852308, 4.46795779229051, 4.54289874938464, 4.69127381231347, 
    4.88911027911278,
  5.31594290645771, 5.00605454456741, 4.79455372505948, 4.68097694456457, 
    4.63086548203189, 4.63211348404195, 4.70096220131872, 4.83925041999867, 
    5.02242318217544,
  5.4455350902829, 5.1479946960376, 4.94692989373408, 4.84147051544417, 
    4.79704625989776, 4.80121777526291, 4.86801953101339, 4.99889544145281, 
    5.16612461065588 ;

 lon_psi =
  -49.8852333380674, -49.4134990783, -48.9252885750958, -48.3992602989844, 
    -47.8355302481014, -47.2493955379091, -46.6658939438917, 
    -46.0892372814687, -45.5120325830865,
  -49.7983157950911, -49.3247798106966, -48.8398016032612, -48.342986239888, 
    -47.8326230768061, -47.2842335118098, -46.7131898670564, 
    -46.1368665842142, -45.5585345385222,
  -49.7053855498322, -49.2347637641474, -48.7584995867321, -48.2911154947519, 
    -47.8255840571535, -47.3132752115364, -46.7583885614251, 
    -46.1855155507126, -45.6087666910297,
  -49.6093094769188, -49.1455616908453, -48.6823286124262, -48.2434477350499, 
    -47.8157175121508, -47.3368626214109, -46.8005639047206, 
    -46.2339656435392, -45.6610892191651,
  -49.5116157313484, -49.0578406650387, -48.6108593350757, -48.1992392899088, 
    -47.8040698339627, -47.3560038362421, -46.8397411992034, 
    -46.2817334429845, -45.7144616601388,
  -49.4130978527148, -48.9715512267185, -48.5432236181582, -48.157749609441, 
    -47.7914291660544, -47.3718463314966, -46.8763887171883, 
    -46.3287048789574, -45.7681251513714,
  -49.3140177675271, -48.8861129495609, -48.4783663090131, -48.1183292012273, 
    -47.7784155436412, -47.3855617349024, -46.9112667193033, 
    -46.3750413836221, -45.8214418668094,
  -49.2140313949058, -48.800251205493, -48.4149755293871, -48.0803543148767, 
    -47.7655736313989, -47.3984121609982, -46.9454778731932, 
    -46.4212551939777, -45.8738023865188,
  -49.1114134802482, -48.7110465771771, -48.3509045159634, -48.042947902838, 
    -47.7534506972285, -47.4120506667142, -46.9808820202716, 
    -46.4686715374539, -45.9246717758002 ;

 lat_u =
  4.50026015768974, 4.0780984466164, 3.68974214127326, 3.40468299651808, 
    3.3129814902132, 3.41691150585875, 3.62519560217182, 3.87989047390449, 
    4.14137956892014,
  4.59238254566534, 4.18045789421623, 3.82366197839628, 3.58064151767931, 
    3.49612877353478, 3.56740723781395, 3.74606091560509, 3.98273132689303, 
    4.23880464487679,
  4.69448024714094, 4.29582982385791, 3.9700878758053, 3.76213646940812, 
    3.68422578107596, 3.72998047498617, 3.88061382432594, 4.09845013231385, 
    4.34722948768657,
  4.80081362351111, 4.41744846877268, 4.11974755822207, 3.93902259705286, 
    3.86689719533252, 3.89459573941108, 4.02122300474378, 4.22095797566988, 
    4.46077875223404,
  4.91028279103098, 4.5434008708195, 4.27045399066847, 4.11102624962995, 
    4.04410176848109, 4.05938233354052, 4.16619703433325, 4.34907154934143, 
    4.57845625173846,
  5.02223425293318, 4.67230453619823, 4.42079265385458, 4.27814193033295, 
    4.21604233174045, 4.22328664371716, 4.31443642590749, 4.48207789365758, 
    4.69972522075001,
  5.13672161055677, 4.80358280192979, 4.57036015808752, 4.44114883552055, 
    4.38372173719402, 4.38636551002045, 4.46576135677245, 4.62004072474511, 
    4.8247714251298,
  5.25503936593683, 4.93779562575485, 4.71981945834291, 4.60153926136824, 
    4.54890641982382, 4.5499233599828, 4.6213529329551, 4.76438643740965, 
    4.95502949463879,
  5.37844473839587, 5.07530405730512, 4.86947605864466, 4.76015859453574, 
    4.71271192334709, 4.7149111507644, 4.78214217754598, 4.91633427367731, 
    5.09175296046628,
  5.52083595106861, 5.22711914551171, 5.02978239041476, 4.92782192147353, 
    4.88703192397131, 4.89456437985436, 4.96239869267397, 5.09088859868507, 
    5.24930495448903 ;

 lon_u =
  -49.9237898688101, -49.4546545157168, -48.96698536448, -48.4275774358079, 
    -47.8351480599858, -47.2309074499535, -46.643036086764, 
    -46.0672576162864, -45.4915757996105,
  -49.842980707126, -49.3697566990597, -48.8824448514824, -48.3707996339772, 
    -47.8346566575698, -47.2673706542632, -46.6895438503016, 
    -46.1126800559703, -45.5345762032174,
  -49.7523350642767, -49.2796997867542, -48.7984554169598, -48.3164422950536, 
    -47.8295409140893, -47.299516062078, -46.7361738159154, 
    -46.1611927695097, -45.5833304453076,
  -49.6576382542949, -49.1900145277432, -48.7198015503493, -48.2668121771525, 
    -47.8209311662385, -47.3256849469602, -46.7798560989976, 
    -46.2097978695312, -45.6347332757956,
  -49.5606015612579, -49.1015053448438, -48.6460520715151, -48.2209564732413, 
    -47.8100630465528, -47.3469200883111, -46.8205065115458, 
    -46.257949189239, -45.687696718153,
  -49.46242589976, -49.0145352399062, -48.5766209132696, -48.1781952646626, 
    -47.7978319205278, -47.3642659584268, -46.8583421884275, 
    -46.3053178009772, -45.7413001098915,
  -49.3636622994392, -48.9288147143841, -48.5105396311338, -48.1378276707736, 
    -47.7849355283593, -47.3788883547697, -46.8939770723734, 
    -46.3519156608304, -45.7948563111196,
  -49.2640882014603, -48.843251893177, -48.4465209608704, -48.0991698335125, 
    -47.7719349395798, -47.3920308130467, -46.928411286042, 
    -46.3981636402373, -45.8478128287319,
  -49.1636901533346, -48.7567993841749, -48.3835003275502, -48.0617952930102, 
    -47.759403574472, -47.4049004685343, -46.9626773290685, 
    -46.4444544908711, -45.8993192181678,
  -49.0551769286559, -48.6607583450266, -48.3157569671346, -48.0231529010941, 
    -47.7477294213616, -47.420507746918, -47.0011296929789, 
    -46.4950092303901, -45.9502684550684 ;

 lat_v =
  4.75220777929874, 4.33368362225529, 3.93117277259219, 3.60396462788413, 
    3.42293421092423, 3.42793878348367, 3.57682549069983, 3.80231802181795, 
    4.0582653916216, 4.31692748101462,
  4.84920710801575, 4.43590445528519, 4.05497458031167, 3.76720838377744, 
    3.61304533984139, 3.60374509448146, 3.71964894896946, 3.92083622959231, 
    4.16417949859427, 4.42223205338393,
  4.94965192436719, 4.5458323096783, 4.1870299316353, 3.9326297619882, 
    3.79939095780102, 3.78057487534026, 3.8700250355361, 4.04813850957202, 
    4.27826988073563, 4.532008476268,
  5.05198586082778, 4.66066069991856, 4.32345025966525, 4.09658208510835, 
    3.97949636614238, 3.95490103797895, 4.02400146123902, 4.18144257367589, 
    4.398046265988, 4.64472633151481,
  5.15568823034591, 4.77900614365996, 4.46219513393646, 4.2578868861457, 
    4.15346173544546, 4.12585398476908, 4.17982997407027, 4.31948909738785, 
    4.52254495098802, 4.75970502494616,
  5.26078645834676, 4.90029796071154, 4.60226052712173, 4.41641799554881, 
    4.3221960128993, 4.29367108700113, 4.3369411174517, 4.46189713901639, 
    4.65162892630642, 4.87691596494309,
  5.36780851194808, 5.02469612606949, 4.74341291332996, 4.57265649933423, 
    4.48695736621102, 4.45924255310396, 4.49565419802866, 4.60907317429049, 
    4.78593272861686, 4.99677389240053,
  5.47810678235593, 5.15342792264811, 4.8862967689691, 4.72774875803058, 
    4.64947387740263, 4.62423610996141, 4.65738860344945, 4.76256655940655, 
    4.92727352848904, 5.12036856633162,
  5.59517589949956, 5.29029794752599, 5.03348295158058, 4.88455414246113, 
    4.81308177445425, 4.79237294745454, 4.82612179262171, 4.92668985027181, 
    5.08041715037122, 5.25065965288912 ;

 lon_v =
  -50.1143422941785, -49.6511435189659, -49.1727309171351, -48.6675090206378, 
    -48.1214396790943, -47.5435905999823, -46.9565038361161, 
    -46.3774472569268, -45.7998879242123, -45.2293070288291,
  -50.0197787930178, -49.5646480096826, -49.083383313994, -48.5926530538427, 
    -48.091194880627, -47.5629485985285, -46.9999954308976, -46.425848099749, 
    -45.8458704738008, -45.282045952558,
  -49.9201627606786, -49.4738617834176, -48.9957594708396, -48.5232950975756, 
    -48.0612469757871, -47.5762000607875, -47.0393611855684, 
    -46.4737759951864, -45.8945143939027, -45.3380383584601,
  -49.8176496612721, -49.3814573760496, -48.9114427180206, -48.4595510252694, 
    -48.0321200802698, -47.5844676435831, -47.0741786843594, 
    -46.5201292760691, -45.9443206426833, -45.3960781461763,
  -49.713465013435, -49.2886682700008, -48.8305312231359, -48.4005762154416, 
    -48.0039362743034, -47.5890503148902, -47.1049468291136, 
    -46.5646547551794, -45.9944819335064, -45.4552482469017,
  -49.6083286186107, -49.195952608216, -48.7525033247034, -48.3453677047605, 
    -47.976696434699, -47.5911192796994, -47.1325107927913, 
    -46.6075300697312, -46.0445094525615, -45.5148795994984,
  -49.502617353849, -49.1031812968281, -48.6764509400914, -48.2929361823008, 
    -47.9503699842966, -47.5917160274988, -47.157900071587, 
    -46.6492476079023, -46.0941207429283, -45.5743318073843,
  -49.3963531065656, -49.0094976700839, -48.6009610718778, -48.2422331189084, 
    -47.9249078593587, -47.5918517504975, -47.182373315302, 
    -46.6906924397669, -46.1432413121865, -45.6328591130416,
  -49.2887503299089, -48.9123695385965, -48.5233262472178, -48.1917300381972, 
    -47.9001414633482, -47.5927194814362, -47.207775772631, 
    -46.7336241824591, -46.1922842813078, -45.6895306741425 ;

 mask_rho =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mask_u =
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mask_v =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mask_psi =
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 angle =
  -0.703507710608412, -0.734199126280519, -0.67352593984004, 
    -0.487320983768581, -0.153817760791567, 0.170849817176119, 
    0.340619724598406, 0.416735450771849, 0.427036372382658, 0.408473084257683,
  -0.747797502777564, -0.717968557937026, -0.633716949282945, 
    -0.445120912447325, -0.156589593857297, 0.126031392236994, 
    0.300671608979915, 0.39008459693982, 0.417744925482352, 0.442546378838024,
  -0.76974843390473, -0.702546165676821, -0.597152289811802, 
    -0.409255142345235, -0.158925711326187, 0.0873955856722987, 
    0.262482494280695, 0.363174063492778, 0.407343232888974, 0.459224015914168,
  -0.78137531191013, -0.688616169295746, -0.566522631409318, 
    -0.381360013438075, -0.160667142931213, 0.0569141373485191, 
    0.229160799607476, 0.338083399983138, 0.395915435621555, 0.466821460696627,
  -0.786560298231328, -0.676197537596091, -0.542029960609056, 
    -0.360449968223552, -0.161778613030964, 0.0338923970995636, 
    0.201411967398258, 0.315423225289811, 0.383256865474535, 0.468242950639523,
  -0.786920000535964, -0.665277079138279, -0.523507383689382, 
    -0.345371991128099, -0.162169505009777, 0.0175098743724356, 
    0.17947396849437, 0.295484637309201, 0.369072384885805, 0.464177238125456,
  -0.7823332062841, -0.655887566864309, -0.510948608436446, 
    -0.335273481296227, -0.161631283151678, 0.00732415720229451, 
    0.163578155379685, 0.278490505905563, 0.352919980202553, 0.454105452457469,
  -0.770262404943912, -0.648231816818805, -0.504919657253734, 
    -0.329837500903909, -0.159742126376036, 0.00358413699336254, 
    0.15425864723804, 0.264755913187296, 0.334121409580397, 0.43516810941705,
  -0.742305905059412, -0.643080583248282, -0.50728404247734, 
    -0.329681702834835, -0.155595916329142, 0.00783567975840999, 
    0.152790250294528, 0.254890560995613, 0.311634053536323, 0.399173394958195,
  -0.653266031694124, -0.643837857657218, -0.524951997135465, 
    -0.33866965838004, -0.146137966573541, 0.0265114531620193, 
    0.163435345267253, 0.250552800732948, 0.282727931115157, 0.304085790441704 ;
}
